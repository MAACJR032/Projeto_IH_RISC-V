`timescale 1ns / 1ps

module Controller (
    //Input
    input halt_reg,
    input logic [6:0] Opcode,
    //7-bit opcode field from the instruction

    //Outputs
    output logic ALUSrc,
    //0: The second ALU operand comes from the second register file output (Read data 2); 
    //1: The second ALU operand is the sign-extended, lower 16 bits of the instruction.
    output logic MemtoReg,
    //0: The value fed to the register Write data input comes from the ALU.
    //1: The value fed to the register Write data input comes from the data memory.
    output logic RegWrite, //The register on the Write register input is written with the value on the Write data input 
    output logic MemRead,  //Data memory contents designated by the address input are put on the Read data output
    output logic MemWrite, //Data memory contents designated by the address input are replaced by the value on the Write data input.
    output logic [1:0] ALUOp,  //00: LW/SW; 01:Branch; 10: R-Type/I-Type 11: JAL/LUI
    output logic Branch,  //0: branch is not taken; 1: branch is taken
    output logic halt
);

  logic [6:0] R_TYPE, I_TYPE, LW, SW, BR, J, JR, HALT;

  assign R_TYPE = 7'b0110011; // add,and,sub,or,xor,slt
  assign I_TYPE = 7'b0010011; // addi,slti,slli,srli,srai
  assign LW = 7'b0000011; // lw
  assign SW = 7'b0100011; // sw
  assign BR = 7'b1100011; // beq,bne,blt,bge
  assign J = 7'b1101111; // jal
  assign JR = 7'b1100111; //jalr
  assign HALT = 7'b0000001; // halt

  assign ALUSrc = (Opcode == LW || Opcode == SW || Opcode == I_TYPE);
  assign MemtoReg = (Opcode == LW);
  assign RegWrite = (Opcode == R_TYPE || Opcode == I_TYPE || Opcode == LW || Opcode == J || Opcode == JR);
  assign MemRead = (Opcode == LW);
  assign MemWrite = (Opcode == SW);
  assign ALUOp[0] = (Opcode == BR || Opcode == J || Opcode == JR);
  assign ALUOp[1] = (Opcode == R_TYPE || Opcode == I_TYPE || Opcode == J || Opcode == JR);
  assign Branch = (Opcode == BR || Opcode == J || Opcode == JR);
  assign halt = (Opcode == HALT) || (halt_reg);

endmodule
